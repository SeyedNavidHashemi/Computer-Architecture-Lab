module or_module(first, second, result);
    input first, second;
    output result;

    assign result = first | second;
endmodule